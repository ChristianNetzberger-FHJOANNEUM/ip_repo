//
// Verilog Module training_lib.circuit_ch1_2e_v
//
// Created:
//          by - net.UNKNOWN (KPERSM7467)
//          at - 10:33:35 03.11.2017
//
// using Mentor Graphics HDL Designer(TM) 2016.2 (Build 5)
//

`resetall
`timescale 1ns/10ps
module circuit_ch1_2e_v ;


// ### Please start your Verilog code here ### 

endmodule
