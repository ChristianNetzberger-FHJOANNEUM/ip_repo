--
-- VHDL Architecture sbus_uart_lib.resync.rtl
--
-- Created:
--          by - net.UNKNOWN (KPERSM7467)
--          at - 11:33:22 08.11.2018
--
-- using Mentor Graphics HDL Designer(TM) 2016.2 (Build 5)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

entity resync is
  port(clk: in std_logic;
       stb_a: in std_logic;
       sync_en: in std_logic;
       stb_s: out std_logic);
end entity resync;

--
architecture rtl of resync is
begin
      
end architecture rtl;

